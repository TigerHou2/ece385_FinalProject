//------------------------------------------------------------------------
//																								--
//			ECE 385 Final Project, Spring 2021										--
//			Tiger Hou																		--
//																								--
//------------------------------------------------------------------------


module FinalProject (

      ///////// Clocks /////////
      input     CLOCK_50,

      ///////// KEY /////////
      input    [ 1: 0]   KEY,

      ///////// SW /////////
      input    [ 9: 0]   SW,

      ///////// LEDR /////////
      output   [ 9: 0]   LEDR,

      ///////// HEX /////////
      output   [ 7: 0]   HEX0,
      output   [ 7: 0]   HEX1,
//      output   [ 7: 0]   HEX2,
      output   [ 7: 0]   HEX3,
      output   [ 7: 0]   HEX4,
//      output   [ 7: 0]   HEX5,

      ///////// SDRAM /////////
      output             DRAM_CLK,
      output             DRAM_CKE,
      output   [12: 0]   DRAM_ADDR,
      output   [ 1: 0]   DRAM_BA,
      inout    [15: 0]   DRAM_DQ,
      output             DRAM_LDQM,
      output             DRAM_UDQM,
      output             DRAM_CS_N,
      output             DRAM_WE_N,
      output             DRAM_CAS_N,
      output             DRAM_RAS_N,

      ///////// VGA /////////
      output             VGA_HS,
      output             VGA_VS,
      output   [ 3: 0]   VGA_R,
      output   [ 3: 0]   VGA_G,
      output   [ 3: 0]   VGA_B,


      ///////// ARDUINO /////////
      inout    [15: 0]   ARDUINO_IO,
      inout              ARDUINO_RESET_N 

);




logic Reset_h, vssig, blank, sync, VGA_Clk;


//=======================================================
//  REG/WIRE declarations
//=======================================================
	logic SPI0_CS_N, SPI0_SCLK, SPI0_MISO, SPI0_MOSI, USB_GPX, USB_IRQ, USB_RST;
	logic [3:0]		hex_num_4, hex_num_3, hex_num_1, hex_num_0; //4 bit input hex digits
	logic [9:0]		drawxsig, drawysig;
	logic [7:0]		Red, Blue, Green;
	logic [15:0]	keycode;
	logic [7:0]		key_p1, key_p2;
	logic [17:0]	P1A, P2A, B1A, B2A;
	logic				P1D, P2D, B1D, B2D;
	logic				BB1, BB2;
	logic	[63:0]	P1C, P2C;
	logic [9:0]		B1X, B1Y, B2X, B2Y;
	logic [9:0]		HP1, HPP1, HP2, HPP2;
	logic [17:0]	addrBG;
	logic				drawBG;

//=======================================================
//  Structural coding
//=======================================================
	assign ARDUINO_IO[10] = SPI0_CS_N;
	assign ARDUINO_IO[13] = SPI0_SCLK;
	assign ARDUINO_IO[11] = SPI0_MOSI;
	assign ARDUINO_IO[12] = 1'bZ;
	assign SPI0_MISO = ARDUINO_IO[12];
	
	assign ARDUINO_IO[9] = 1'bZ; 
	assign USB_IRQ = ARDUINO_IO[9];
		
	//Assignments specific to Circuits At Home UHS_20
	assign ARDUINO_RESET_N = USB_RST;
	assign ARDUINO_IO[7] = USB_RST;//USB reset 
	assign ARDUINO_IO[8] = 1'bZ; //this is GPX (set to input)
	assign USB_GPX = 1'b0;//GPX is not needed for standard USB host - set to 0 to prevent interrupt
	
	//Assign uSD CS to '1' to prevent uSD card from interfering with USB Host (if uSD card is plugged in)
	assign ARDUINO_IO[6] = 1'b1;
	
	//HEX drivers to convert numbers to HEX output
	HexDriver hex_driver4 (hex_num_4, HEX4[6:0]);
	assign HEX4[7] = 1'b1;
	
	HexDriver hex_driver3 (hex_num_3, HEX3[6:0]);
	assign HEX3[7] = 1'b1;
	
	HexDriver hex_driver1 (hex_num_1, HEX1[6:0]);
	assign HEX1[7] = 1'b1;
	
	HexDriver hex_driver0 (hex_num_0, HEX0[6:0]);
	assign HEX0[7] = 1'b1;
	
	
	//Assign one button to reset
	assign {Reset_h}=~ (KEY[0]);

	//Our A/D converter is only 12 bit
	assign VGA_R = Red[7:4];
	assign VGA_B = Blue[7:4];
	assign VGA_G = Green[7:4];
	
	// Terrain data assignments
	logic [479:0]	T1O, T2O, terrain_out;
	logic [9:0]		terrain_addr;
	logic [9:0]		terrain_height;
	logic [17:0]	addrTerrain;
	logic				drawTerrain;
	
	always_ff @ (negedge CLOCK_50)
	begin
		terrain_addr <= drawxsig - 1'b1;
	end
	
	// Player keycode assignments
	assign key_p1 = keycode[15:8];
	assign key_p2 = keycode[7:0];
	
	// Player controls
	assign P1C = {8'd26, 8'd22, 8'd04, 8'd07, 8'd20, 8'd08, 8'd30, 8'd32}; // W,S,A,D,Q,E,1,3
	assign P2C = {8'd12, 8'd14, 8'd13, 8'd15, 8'd24, 8'd18, 8'd37, 8'd38}; // I,K,J,L,U,O,8,9
	
	// Scoring
	logic				drawScore;
	logic [17:0]	addrScore;
	
	// Debug
	assign LEDR = HPP1;
	
	
	finalsoc u0 (
		.clk_50_clk                        (CLOCK_50),  		//clk_50.clk
		.reset_50_reset_n                  (1'b1),         	//reset_50.reset_n
		.altpll_0_locked_conduit_export    (),						//altpll_0_locked_conduit.export
		.altpll_0_phasedone_conduit_export (),						//altpll_0_phasedone_conduit.export
		.altpll_0_areset_conduit_export    (),						//altpll_0_areset_conduit.export
		.key_external_connection_export    (KEY),					//key_external_connection.export

		//SDRAM
		.sdram_clk_clk(DRAM_CLK),										//clk_sdram.clk
		.sdram_wire_addr(DRAM_ADDR),									//sdram_wire.addr
		.sdram_wire_ba(DRAM_BA),										//.ba
		.sdram_wire_cas_n(DRAM_CAS_N),								//.cas_n
		.sdram_wire_cke(DRAM_CKE),										//.cke
		.sdram_wire_cs_n(DRAM_CS_N),									//.cs_n
		.sdram_wire_dq(DRAM_DQ),										//.dq
		.sdram_wire_dqm({DRAM_UDQM,DRAM_LDQM}),					//.dqm
		.sdram_wire_ras_n(DRAM_RAS_N),								//.ras_n
		.sdram_wire_we_n(DRAM_WE_N),									//.we_n

		//USB SPI	
		.spi0_SS_n(SPI0_CS_N),
		.spi0_MOSI(SPI0_MOSI),
		.spi0_MISO(SPI0_MISO),
		.spi0_SCLK(SPI0_SCLK),
		
		//USB GPIO
		.usb_rst_export(USB_RST),
		.usb_irq_export(USB_IRQ),
		.usb_gpx_export(USB_GPX),
		
		//LEDs and HEX
		.hex_digits_export({hex_num_4, hex_num_3, hex_num_1, hex_num_0}),
//		.leds_export({hundreds, signs, LEDR}),
		.keycode_export(keycode)
		
	 );


//instantiate a vga_controller, ball, and color_mapper here with the ports.

player P1				(	.clk(CLOCK_50), .reset(Reset_h), .frame_clk(VGA_VS), .terrain_data(terrain_out),
								.keycode(key_p1), .DrawX(drawxsig), .DrawY(drawysig), .ID(1'b0), .controls(P1C),
								.DX(B2X), .DY(B2Y), .Dboomed(BB2), .BX(B1X), .BY(B1Y), .boomed(BB1), .HP(HP1), .HPP(HPP1),
								.drawPlayer(P1D), .drawBomb(B1D), .addrPlayer(P1A), .addrBomb(B1A),
								.terrain_out(T1O));
								
player P2				(	.clk(CLOCK_50), .reset(Reset_h), .frame_clk(VGA_VS), .terrain_data(terrain_out),
								.keycode(key_p2), .DrawX(drawxsig), .DrawY(drawysig), .ID(1'b1), .controls(P2C),
								.DX(B1X), .DY(B1Y), .Dboomed(BB1), .BX(B2X), .BY(B2Y), .boomed(BB2), .HP(HP2), .HPP(HPP2),
								.drawPlayer(P2D), .drawBomb(B2D), .addrPlayer(P2A), .addrBomb(B2A),
								.terrain_out(T2O));
				
vga_controller VGA	(	.Clk(CLOCK_50), .Reset(Reset_h), .hs(VGA_HS), .vs(VGA_VS),
								.pixel_clk(VGA_Clk), .blank, .sync, .DrawX(drawxsig), .DrawY(drawysig)  );

color_mapper CMAP		(	.clk(CLOCK_50), 
								.P1A, .P2A, .B1A, .B2A, .addrBG, .addrTerrain, .addrScore,
								.P1D, .P2D, .B1D, .B2D, .drawBG, .drawTerrain, .drawScore,
								.blank, .Red, .Green, .Blue  );

terrain TERRAIN		(	.clk(CLOCK_50), .we((~B1D)&(~B2D)&blank), .reset(Reset_h), 
								.DrawX(drawxsig), .DrawY(drawysig), .terrain_in(T1O&T2O), 
								.read_addr(drawxsig), .write_addr(terrain_addr), .rngSeed(SW), 
								.terrain_out, .terrain_height, .addrTerrain, .drawTerrain);

background BACKGROUND(	.mapSelect(SW[9]), .DrawX(drawxsig), .DrawY(drawysig), .drawBG, .addrBG);

scoreboard SCOREBOARD(	.DrawX(drawxsig), .DrawY(drawysig), .HP1, .HPP1, .HP2, .HPP2, .drawScore, .addrScore);

endmodule
